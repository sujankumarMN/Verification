package mul_package;

	class mul_transaction;
		bit [1:0]A;
		bit [1:0]B;
		bit [3:0]product;
		bit loadA,loadB,decB,loadF,clear,zero,start;
		bit [1:0]P;
		bit [1:0]Q;
	endclass
endpackage
